`FOO

`define BAR 666
`BAR

`undefineall

`ifdef FOO

123
`BAR

`endif
