package pkg;

localparam FOO = 1;

endpackage