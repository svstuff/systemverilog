function foo;
   a.b[i][j] = c[i][8*j +:8];
endfunction
