function int clazz::func(string name);
   !this.foo();
endfunction
