`define SIZE 42
`define D(a) `SIZE``a
`D('d0)
