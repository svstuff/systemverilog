function int clazz::func(string name);
  // call static function 'func' in class 'clazz' in package 'pkg'
  pkg::clazz::func();
endfunction
