`define append(a,b) a``b
`append(foo,bar)
