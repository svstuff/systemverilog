/** **/
