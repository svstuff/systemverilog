`define DEF(A,B,C) a_``B_``C

`DEF(a, b, c)
