function int func;
   --yo;
endfunction
