typedef mailbox #(foo_t) bar_t;
