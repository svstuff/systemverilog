`define DEF1(A,B) `DEF2(B,A)
`define DEF2(A,B) A+B

`DEF1(a,b)
