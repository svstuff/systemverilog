function void func();
      foo = 64'(bar[0]);
endfunction
