// single line comment with no newline