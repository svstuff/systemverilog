module adder2(a, b, c);
endmodule
