`define DEF1(A,B) A `DEF2(1+B)
`define DEF2(C) (C)

`DEF1(a,b)
