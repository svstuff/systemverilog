function void connect_phase;
  reg2apb_adapter reg2apb = new;
endfunction
