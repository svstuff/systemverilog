function int clazz::func(string name);
   this.randomize(this.foo);
   void'(this.jcb_rq.deep_copy(jcb_rq_copy));
endfunction
