module mod1 ();
endmodule : label1

module mod2 (a,b,c) ;
endmodule
