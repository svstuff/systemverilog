`define FOO $display("yo")

`FOO(foo)
