
// This test does nothing but include uvm macros.
`include "uvm_macros.svh"
