function void clazz::func();

  arg = { arg, string'(char) };

endfunction
