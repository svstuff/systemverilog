`define YO

foo `YO bar
