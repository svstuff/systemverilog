function foo;
   if( !bar() ) return;
endfunction
