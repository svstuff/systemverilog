`define FOO(a,b) a + b
`FOO( {0,1,2}, 42 )