
function foo;
   symbol = {symbol[6:0], rx};
endfunction
