`define UVM_NAME UVM
`define UVM_MAJOR_REV 1
`define UVM_MINOR_REV 1
`define UVM_FIX_REV d

`define UVM_VERSION_STRING `"`UVM_NAME``-```UVM_MAJOR_REV``.```UVM_MINOR_REV`UVM_FIX_REV`"

`UVM_VERSION_STRING
