`define BAR 64
`define FOO(V) `BAR``V

`FOO('d0)
