class class_name extends base_name;

  extern function void foo(pkg1::typ1 a, output pkg2::typ2 b[pkg3::typ3]);

endclass
