`define FOO(a,b) \
"This is \"line\" ..." a\
"and this \"is\" line ..." b

`FOO(2,3)