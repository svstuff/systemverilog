`define FOO(a) a+a+ a+ a +a +!a+a!+ab+ba+bab+_a+a_+a1+1a
`FOO(c)
