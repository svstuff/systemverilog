function void clazz::func(ref string param[string]);
endfunction

function logic [15:0] myfunc2;
  input int x;
  input int y;
endfunction

function [3:0][7:0] myfunc4(input [3:0][7:0] a, b[3:0]);

endfunction
