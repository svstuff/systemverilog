
`define FOO(TYPE,ARG,FLAG) `M_UVM_``TYPE(ARG,FLAG)
`define M_UVM_ARRAY(arg1, arg2) yo

`FOO(ARRAY, byte_valid, UVM_NOPACK)
