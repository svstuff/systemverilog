function int func();
  void'(std::randomize(yo));
endfunction
