`define YO veryverylongnamesothatsubsequenttokenswouldgetthewrongcolumn
`YO 1 `YO