function int clazz::func(string name);
  foo(data[7:0]);
endfunction
