`define FOO(a,b) a + b
`define BAR(c) [c]
`FOO(foo,`BAR(bar))