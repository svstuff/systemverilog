`define YO(a,b,c) a + b + c
`YO(foo,bar,yo)