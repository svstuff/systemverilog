`define D(a) /*foo a bar*/ a b c
`D(42)