class clazz #(type T = data);
endclass
