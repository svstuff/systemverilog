`define FOO(yo) yo + `BAR(bar)
`define BAR(yo) yo
`FOO(foo)