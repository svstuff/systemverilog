class test;
  virtual function bit test();
      return (randomize(null));
  endfunction
endclass
