import "DPI-C" function int system(string  s);
