task foo();
  pkg::clazz1#(42)::method1().method2().method3();
//  pkg::clazz1#(42)::clazz2::staticmethod().method1().method2().member1.member2
endtask
