module test();
input wire [WIDTH-1:0]  array_with_unpacked_dimension [0:SOMENUM-1];
endmodule
