function foo;
   // note: a[0].b is an expression / hierarchical-id.
   // [i] is the loop variable part of the foreach.
   foreach ( a[0].b[i] )
     begin
     end
endfunction
