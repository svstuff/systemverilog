function int clazz::func(string name);
endfunction
