`define BAR(a) f(a) f(a,x) f(x,a) f(x,a,y)
`BAR(c)
