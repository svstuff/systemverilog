task test();
  foreach (testarray[i]) begin
  end
endtask : test
