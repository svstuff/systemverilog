function int clazz::func(string name);
   this.randomize(this.foo);
endfunction
