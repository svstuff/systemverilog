`define append(a,b) ab a``b+a+b
`append(foo,bar)
