function void clazz::func(ref string param[string]);
endfunction
