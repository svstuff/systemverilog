?
!
!=
!==
!=?
%
&
&&
*
**
+
++
-
--
->
/
<
<->
<<
<<<
<=
==
===
==?
>
>=
>>
>>>
^
^~
| 
||
~
~&
~^
~|
=
+=
-=
*=
/=
%=
&=
|=
^=
<<=
>>=
<<<=
>>>=
