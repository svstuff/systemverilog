
function foo;
   a.b.c = 0;
endfunction
