`define FOO( a, b=c(d,e) ) a+b
`FOO(1,)
