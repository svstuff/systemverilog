æøå this shouldn't be included!