
function foo;
   a = 0
endfunction
