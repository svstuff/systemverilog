typedef uvm_component_registry #(producer #(T),"producer #(T)") type_id;
