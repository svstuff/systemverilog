
localparam FOO = BAR >>> 1;
localparam FOO = BAR <<< 1;
