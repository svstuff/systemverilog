`define FOO(a,b) a + b
`define BAR(c) [c]
`define YO(d) {d}
`FOO(foo,`BAR(`YO(bar)))