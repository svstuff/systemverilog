/* multiline comment */