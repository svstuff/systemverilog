task clazz::func(string name);
  if (env[i].name == name)
    return ;
endtask
