package pkg;

clazz#(param1,param2) myvar;
   
endpackage
