`define FOO( a=1, b=2 ) a+b
`FOO(,)
