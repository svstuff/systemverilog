`define D(a,b) a+b
`D(1 /* comment */, 2)
