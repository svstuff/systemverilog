function int func();
  q = test.find_first_index with (item.A == test2.B);
endfunction
