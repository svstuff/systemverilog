interface vpe_ace4_lite_slave_if (input bit FOO, input bit BAR);

endinterface
