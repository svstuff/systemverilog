`define YO(a,b) a + b
`YO(foo,bar)