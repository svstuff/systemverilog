task clazz::func();
  if ( a.randomize() with {} ) begin
  end
endtask
