`ifdef FOO
  foo(" ")
`endif
bar
