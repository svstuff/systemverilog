function void build_phase();
  uvm_config_db#(apb_vif)::get();
endfunction
