task clazz::func(string name);
  foreach (env[i])
    if (env[i] == name)
      return ;
endtask
