function int clazz::func(string name);
   if ( !this.randomize(this.foo) ) bar();
endfunction
