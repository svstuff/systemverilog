some
tokens
here