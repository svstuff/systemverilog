function int clazz::func();
  string parts[$];
endfunction
