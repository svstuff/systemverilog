function void clazz::func();

  if( max_severity inside { c, d } && e == (f + g + 1) )
    return;

endfunction
