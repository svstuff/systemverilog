`define FOO(a,b) [a]+[b]
`FOO( "abc,\"def\"", 2 )