task clazz;
  int foo[ bar ] =
    '{
       YO  : 3
     };
endtask
