function int func();
  bar().zoo();
endfunction
