`define DEF1 `DEF2 bar
`define DEF2 foo

`DEF1
