function int clazz::func(string name);
  foreach ( events[event_index] ) begin
    -> events[event_index];
  end
endfunction
