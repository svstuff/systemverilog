/********/
/* multiline comment */
/********/
