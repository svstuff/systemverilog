function foo;
   foreach ( a.b[i,j] )
     begin
     end
endfunction
