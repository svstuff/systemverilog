function foo;
  yo = new this;
endfunction
