`define DEF1(A) `DEF2(A) B
`define DEF2(B) B
`define A yo

`DEF1(`A)
