`ifdef FOO

`FOO

`undef FOO

`ifdef FOO
123
`endif

`endif
