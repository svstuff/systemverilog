single_line_comment // some line comment
end_of_single_line_comment

simple_comment /* comment */ end_of_simple_comment

simple_comment_2 /* comment * / */ end_of_simple_comment_2

multi_line_comment /* comment line 1
comment line 2
comment line 3 */ end_of_multi_line_comment
