class Foo extends pkg::Bar;

endclass // Foo
