function int clazz::func(string name);
  clazz::member.size();
endfunction
