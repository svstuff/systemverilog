function void func();
   // Casting
   foo = 64'(bar[0]);
endfunction
