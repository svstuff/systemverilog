function int func();
  void'(std::randomize(yo));
  void'( randomize() );
endfunction
