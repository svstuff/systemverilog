3'h3:// 8 bits
1:/2
1:// comment
1:/* comment */
