`define D(a,b) a+b
`D(1 /* comment , with a comma */, 2)

