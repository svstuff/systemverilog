function int clazz::func(string name);
  super.new(name);
endfunction
