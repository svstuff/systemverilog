
function foo;
   a = b[i]++;
endfunction
