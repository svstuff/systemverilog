function int clazz::func(string name);
  return (yo++);
endfunction
