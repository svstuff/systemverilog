`ifdef FOO

`BAR

`endif
