
function foo;
   env[i].memb = 0;
endfunction
