typedef struct {
  foo_t foo;
  longint unsigned bar;
} yo_t;
