`define D(a) "foo a bar"+a
`D(42)