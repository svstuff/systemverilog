function int func();
  std::randomize(yo);
endfunction
