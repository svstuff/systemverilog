function int clazz::func(string name);
  foreach (foo[0][b]) return;
endfunction
