`define D(b) a b c // foo b bar
`D(42)