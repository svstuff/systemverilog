virtual class lower extends uvm_component implements yoyo_uvm_sucks;
  function new (string name, uvm_component parent);
    super.new(name, parent);
  endfunction
endclass

module top;
  initial begin
  end
endmodule
