
function foo;
   m_isr [ TX_ISR ] = 0;
endfunction
