`include "uvm_macros.svh"

    `M_UVM_FIELD_QDA_INT(ARRAY, byte_valid,      UVM_DEFAULT|UVM_NOCOMPARE|UVM_NOPACK)
