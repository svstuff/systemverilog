`define YO(a)

foo `YO(1) bar
